`timescale 1ns/1ns       // Задаёт единицы времени симуляции: 1 нс шаг моделирования

`define clk_period 20    // Определяет период тактового сигнала (20 нс = 50 МГц)

module key_led_top_tb;   // Тестбенч для верхнего уровня key_led_top

	//------------------------------------------------------------
	// Объявление сигналов тестовой среды
	//------------------------------------------------------------
	reg Clk;              // тактовый сигнал 50 МГц
	reg Rst_n;            // активный низкий сброс
	
	wire key_in0;         // сигнал первой кнопки
	wire key_in1;         // сигнал второй кнопки
	reg press0, press1;   // управляющие сигналы для моделей кнопок (эмулируют нажатие)
	
	wire [1:0] led;       // выходные светодиоды

	//------------------------------------------------------------
	// Инстанцирование тестируемого модуля (DUT)
	//------------------------------------------------------------
	key_led_top key_led_top0(
		.Clk(Clk),
		.Rst_n(Rst_n),
		.key_in0(key_in0),
		.key_in1(key_in1),
		.led(led)
	);
	
	//------------------------------------------------------------
	// Модели кнопок — эмулируют дребезг при нажатии
	//------------------------------------------------------------
	key_model key_model0(
		.press(press0),    // внешний управляющий сигнал из тестбенча
		.key(key_in0)      // выход дребезжащего сигнала на вход FPGA
	);
	
	key_model key_model1(
		.press(press1),
		.key(key_in1)
	);
	
	//------------------------------------------------------------
	// Генератор системного тактового сигнала
	//------------------------------------------------------------
	initial Clk = 1;
	always #(`clk_period/2) Clk = ~Clk;  // генерация 50 МГц (20 нс период)

	//------------------------------------------------------------
	// Последовательность теста
	//------------------------------------------------------------
	initial begin
		// 1️⃣ Начальное состояние
		Rst_n  = 1'b0;   // активируем сброс
		press0 = 0;      // кнопки не нажаты
		press1 = 0;
		
		// 2️⃣ Ждём немного, потом снимаем сброс
		#(`clk_period*10)
		Rst_n = 1'b1;
		#(`clk_period*10 + 1);	
		
		// 3️⃣ Первое нажатие кнопки 0 (увеличить счётчик)
		press0 = 1;                    // активируем кнопку
		#(`clk_period*3)
		press0 = 0;                    // отпускаем
		#80_000_000;                   // ждём 80 мс (симулируем задержку пользователя)
		
		// 4️⃣ Второе нажатие кнопки 0
		press0 = 1;
		#(`clk_period*3)
		press0 = 0;
		#80_000_000;
		
		// 5️⃣ Первое нажатие кнопки 1 (уменьшить счётчик)
		press1 = 1;
		#(`clk_period*3)
		press1 = 0;
		#80_000_000;
		
		// 6️⃣ Второе нажатие кнопки 1
		press1 = 1;
		#(`clk_period*3)
		press1 = 0;
		#80_000_000;
		
		// 7️⃣ Остановка симуляции
		$stop;		
	end

endmodule
