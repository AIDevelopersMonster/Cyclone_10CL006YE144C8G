
//====================================================
// Название модуля: key_led_top
// Назначение: Верхний уровень проекта — обработка нажатий кнопок
//              (фильтрация дребезга) и управление светодиодами
// Автор: (твой авторский блок)
// Версия: 1.0
// Дата: (укажи дату)
//====================================================
module key_led_top(
    Clk,     // вход системного тактового сигнала (50 МГц)
    Rst_n,   // системный сброс (активный низкий уровень)
    key_in0, // вход кнопки S0
    key_in1, // вход кнопки S1
    led      // выход на два светодиода
);

    //------------------------------------------------
    // Объявление входов и выходов
    //------------------------------------------------
    input Clk;          // системный тактовый сигнал
    input Rst_n;        // сигнал сброса (активный 0)
    input key_in0;      // кнопка 0
    input key_in1;      // кнопка 1
    output [1:0] led;   // два светодиода

    //------------------------------------------------
    // Промежуточные сигналы
    //------------------------------------------------
    wire key_flag0, key_flag1;   // флаги события нажатия/отпускания кнопки
    wire key_state0, key_state1; // текущее стабильное состояние кнопки

    //------------------------------------------------
    // Подключение фильтра дребезга для кнопки 0
    //------------------------------------------------
    key_filter key_filter0(
        .Clk(Clk),            // системный такт
        .Rst_n(Rst_n),        // сброс
        .key_in(key_in0),     // вход кнопки
        .key_flag(key_flag0), // выход флага события
        .key_state(key_state0)// выход состояния кнопки
    );

    //------------------------------------------------
    // Подключение фильтра дребезга для кнопки 1
    //------------------------------------------------
    key_filter key_filter1(
        .Clk(Clk),
        .Rst_n(Rst_n),
        .key_in(key_in1),
        .key_flag(key_flag1),
        .key_state(key_state1)
    );

    //------------------------------------------------
    // Подключение контроллера светодиодов
    // Он получает обработанные сигналы кнопок
    // и формирует сигналы на выводы светодиодов.
    //------------------------------------------------
    led_ctrl led_ctrl0(
        .Clk(Clk),              // системный такт
        .Rst_n(Rst_n),          // сброс
        .key_flag0(key_flag0),  // флаг кнопки 0
        .key_flag1(key_flag1),  // флаг кнопки 1
        .key_state0(key_state0),// состояние кнопки 0
        .key_state1(key_state1),// состояние кнопки 1
        .led(led)               // выход на светодиоды
    );

endmodule
