`timescale 1ns/1ns   // 1 нс — единица времени симуляции

//------------------------------------------------------------
// Модель кнопки с дребезгом
// Используется в тестбенче для проверки фильтрации
//------------------------------------------------------------
module key_model(
	input  press,  // сигнал "нажать кнопку" из тестбенча
	output reg key // выход "реального" сигнала кнопки (с дребезгом)
);
	
	reg [15:0] myrand; // переменная для случайной задержки дребезга
	
	//------------------------------------------------------------
	// Инициализация — кнопка по умолчанию не нажата
	//------------------------------------------------------------
	initial begin
		key = 1'b1; // уровень 1 = кнопка отпущена
	end
    
	//------------------------------------------------------------
	// Реакция на нажатие сигнала press
	// При каждом фронте вверх выполняется задача press_key
	//------------------------------------------------------------
	always@(posedge press)
		press_key;

	//------------------------------------------------------------
	// Задача моделирования нажатия с дребезгом
	//------------------------------------------------------------
	task press_key;
		begin
			//----------------------------------------------------
			// Этап 1. Симуляция дребезга при нажатии
			//----------------------------------------------------
			repeat(50) begin
				myrand = {$random} % 65536;  // случайная задержка (0–65535 нс)
				#myrand key = ~key;          // инверсия сигнала (имитация дребезга)
			end
			
			key = 0;          // после дребезга кнопка "нажата"
			#25_000_000;      // удержание кнопки ~25 мс
			
			//----------------------------------------------------
			// Этап 2. Симуляция дребезга при отпускании
			//----------------------------------------------------
			repeat(50) begin
				myrand = {$random} % 65536;
				#myrand key = ~key;
			end
			
			key = 1;          // кнопка "отпущена"
			#25_000_000;      // пауза перед возможным следующим нажатием
		end	
	endtask

endmodule
