`timescale 1ns/1ns      // Задает единицы времени и шаг симуляции
                        // 1 нс = базовая единица, шаг моделирования = 1 нс

`define clk_period 20   // Константа: период тактового сигнала = 20 нс (50 МГц)

module key_filter_tb;   // Тестбенч для проверки модуля key_filter

	//------------------------------------------------------------
	// Объявление тестовых сигналов
	//------------------------------------------------------------
	reg Clk;             // системный тактовый сигнал
	reg Rst_n;           // сигнал сброса (активный низкий)
	wire key_in;         // вход от кнопки (будет приходить из модели)
	// reg key_in;        // можно было бы вручную управлять без модели

	wire key_flag;       // выходной флаг события (нажатие/отпускание)
	wire key_state;      // текущее состояние кнопки (0 — нажата, 1 — отпущена)

	//------------------------------------------------------------
	// Подключаем тестируемый модуль (Device Under Test)
	//------------------------------------------------------------
	key_filter key_filter0(
		.Clk(Clk),
		.Rst_n(Rst_n),
		.key_in(key_in),
		.key_flag(key_flag),
		.key_state(key_state)
	);
	
	//------------------------------------------------------------
	// Подключаем модель кнопки
	// Она создаёт дребезг при каждом нажатии
	//------------------------------------------------------------
	key_model key_model(
		.key(key_in)      // выход модели подключен к входу фильтра
	);
	
	//------------------------------------------------------------
	// Генератор системного такта (50 МГц)
	//------------------------------------------------------------
	initial Clk = 1;
	always #(`clk_period/2) Clk = ~Clk;

	//------------------------------------------------------------
	// Последовательность теста
	//------------------------------------------------------------
	initial begin
		Rst_n = 1'b0;                       // активируем сброс
		#(`clk_period * 10) Rst_n = 1'b1;   // снимаем сброс после 10 тактов
		#(`clk_period * 10 + 1);            // подождём немного
	end

endmodule
